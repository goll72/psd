library work;

package attrs is
    constant CPU_N_BITS : natural := 8;
end package;
