package morse_attrs is
    constant COUNTER_CLK_BITS : integer := 26;
    constant MORSE_MAX_LEN : integer := 11;
    constant MORSE_MAX_LEN_BITS : integer := 4;
end package;
