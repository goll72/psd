package morse_attrs is
    -- synthesis translate_off
    constant COUNTER_CLK_BITS : integer := 3;
    -- synthesis translate_on
    -- synthesis read_comments_as_hdl on
    -- constant COUNTER_CLK_BITS : integer := 25;
    -- synthesis read_comments_as_hdl off
    constant MORSE_MAX_LEN : integer := 4;
    constant MORSE_MAX_LEN_BITS : integer := 3;
end package;
